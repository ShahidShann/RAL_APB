package apb_pkg;
   
`include "uvm_macros.svh" 
 import uvm_pkg::*;
 import ral_pkg::*;
 import agent2_pkg::*;
 import pas_agent_pkg::*;

  `include "apb_seq_item.sv"
  `include "adapter.sv"
  `include "apb_driver.sv"
  `include "apb_monitor.sv"
  `include "apb_sequencer.sv"
  `include "apb_agent.sv"
  `include "scoreboard.sv"
  `include "env.sv"
  `include "apb_base_seq.sv"
  `include "apb_rst_seq.sv"
  `include "apb_reg_seq.sv"

  
  
endpackage
