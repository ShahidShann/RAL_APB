package agent2_pkg;
   
`include "uvm_macros.svh" 
 import uvm_pkg::*;
 import ral_pkg::*;

 `include "seq_item.sv" 
 `include "driver.sv"
 `include "monitor.sv"
 `include "agent.sv"
 `include "seq.sv"
endpackage
