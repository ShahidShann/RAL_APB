package test_pkg;
   
`include "uvm_macros.svh" 
 import uvm_pkg::*;
 import ral_pkg::*;
 //`include "scoreboard.sv"
 import apb_pkg::*;
 import agent2_pkg::*;

 `include "apb_base_test.sv"
 `include "apb_test1.sv"
 `include "apb_test2.sv"
  
endpackage
