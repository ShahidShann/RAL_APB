package pas_agent_pkg;
   
`include "uvm_macros.svh" 
 import uvm_pkg::*;
 import ral_pkg::*;
 import agent2_pkg::*;

 `include "pas_monitor.sv"
 `include "pas_agent.sv"
endpackage
